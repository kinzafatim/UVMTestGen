```systemverilog
package tb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "interface.sv"
  `include "and_sequence_item.sv"
  `include "and_sequence.sv"
  `include "and_sequencer.sv"
  `include "and_driver.sv"
  `include "and_monitor.sv"
  `include "and_agent.sv"
  `include "and_env.sv"
  `include "and_scoreboard.sv"
  `include "and_coverage.sv"
  `include "and_test.sv"

endpackage
```